`timescale 1ns / 1ps
//-----------------------------------------------------------------------
//	File:		$RCSfile: Timer.V,v $
//	Version:	$Revision: 1.0 $
//	Desc:		A basic timer module
//	Author:		Farzad Fatollahi-Fard
//	Copyright:	Copyright 2008 UC Berkeley
//	This copyright header must appear in all derivative works.
//-----------------------------------------------------------------------


//-----------------------------------------------------------------------
//	Module:		Timer
//	Desc:		A Timer that counts down from a given input
//	Ex:		T Minus 10, 9, 8, 7, 6, ...
//-----------------------------------------------------------------------
module Timer(Clock, In, Out);
	//---------------------------------------------------------------
	//	I/O
	//---------------------------------------------------------------
	input Clock;
	input [31:0] In;
	output reg Out;
	//---------------------------------------------------------------
	 
	//---------------------------------------------------------------
	//	Regs
	//---------------------------------------------------------------
	reg [31:0] Current;
	//---------------------------------------------------------------

	//---------------------------------------------------------------
	//	Behavioral Timer
	//---------------------------------------------------------------
	always @ (posedge Clock) begin
		Current = (Current != 32'b0) ? (Current - 1) : 32'b0;
		Out = (Current == 32'b0) ? 1'b1 : 1'b0;
	end
	 
	always @ (In) begin
		Current = In;
		Out = 1'b0;
	end
	//---------------------------------------------------------------

endmodule
//-----------------------------------------------------------------------
